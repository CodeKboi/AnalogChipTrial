magic
tech sky130A
magscale 1 2
timestamp 1740587512
<< nwell >>
rect 1128 -216 1180 -214
<< pwell >>
rect 1646 -1362 1698 -1360
rect 1568 -1722 1746 -1686
<< psubdiff >>
rect 1568 -1722 1746 -1686
<< viali >>
rect 1388 -582 1440 -170
rect 1078 -1732 1222 -1682
rect 1568 -1722 1746 -1686
rect 694 -2080 1150 -2042
rect 1800 -2084 2256 -2046
rect 594 -2438 2508 -2358
<< metal1 >>
rect 1324 184 1524 384
rect 1378 -102 1458 184
rect 1632 -100 1708 -96
rect 1124 -104 1292 -102
rect 1116 -148 1292 -104
rect 1376 -148 1458 -102
rect 1116 -186 1192 -148
rect 1376 -170 1456 -148
rect 1534 -152 1708 -100
rect 1116 -214 1230 -186
rect 1376 -198 1388 -170
rect 1116 -296 1128 -214
rect 1118 -550 1128 -296
rect 1108 -580 1128 -550
rect 1182 -580 1230 -214
rect 1282 -578 1388 -198
rect 1108 -600 1230 -580
rect 1376 -582 1388 -578
rect 1440 -198 1456 -170
rect 1440 -578 1544 -198
rect 1632 -210 1708 -152
rect 1600 -228 1714 -210
rect 1600 -576 1650 -228
rect 1706 -576 1714 -228
rect 1440 -582 1456 -578
rect 1108 -632 1184 -600
rect 1108 -682 1286 -632
rect 1118 -684 1286 -682
rect 1376 -686 1456 -582
rect 1600 -586 1714 -576
rect 1638 -634 1714 -586
rect 1540 -678 1714 -634
rect 1540 -686 1708 -678
rect 736 -1266 1278 -1260
rect 1880 -1262 2084 -1258
rect 730 -1312 1278 -1266
rect 730 -1580 934 -1312
rect 1318 -1344 1490 -1268
rect 1530 -1314 2084 -1262
rect 1094 -1354 1196 -1352
rect 1094 -1374 1220 -1354
rect 1094 -1528 1112 -1374
rect 1168 -1528 1220 -1374
rect 1094 -1542 1220 -1528
rect 1142 -1544 1220 -1542
rect 1272 -1552 1538 -1344
rect 1588 -1348 1700 -1344
rect 1588 -1360 1702 -1348
rect 1588 -1532 1646 -1360
rect 1698 -1532 1702 -1360
rect 1588 -1546 1702 -1532
rect 1588 -1548 1700 -1546
rect 1878 -1548 2084 -1314
rect 730 -1632 1272 -1580
rect 948 -1682 1232 -1666
rect 948 -1732 1078 -1682
rect 1222 -1732 1232 -1682
rect 948 -1748 1232 -1732
rect 440 -1902 534 -1894
rect 440 -1962 456 -1902
rect 518 -1962 534 -1902
rect 440 -1970 534 -1962
rect 458 -2272 502 -1970
rect 961 -2015 1043 -1748
rect 569 -2042 1223 -2015
rect 569 -2080 694 -2042
rect 1150 -2080 1223 -2042
rect 569 -2097 1223 -2080
rect 1318 -2126 1490 -1552
rect 1880 -1576 2084 -1548
rect 1698 -1580 2084 -1576
rect 1538 -1606 2084 -1580
rect 1538 -1628 2080 -1606
rect 1532 -1686 1834 -1672
rect 1532 -1722 1568 -1686
rect 1746 -1722 1834 -1686
rect 1532 -1738 1834 -1722
rect 1768 -2031 1834 -1738
rect 2546 -1886 2646 -1878
rect 2546 -1896 2574 -1886
rect 2546 -1954 2568 -1896
rect 2546 -1964 2574 -1954
rect 2626 -1964 2646 -1886
rect 2546 -1968 2646 -1964
rect 1571 -2046 2373 -2031
rect 1571 -2084 1800 -2046
rect 2256 -2084 2373 -2046
rect 1571 -2097 2373 -2084
rect 544 -2214 2534 -2126
rect 1318 -2216 1490 -2214
rect 548 -2358 2538 -2266
rect 2574 -2268 2618 -1968
rect 548 -2438 594 -2358
rect 2508 -2438 2538 -2358
rect 548 -2498 2538 -2438
rect 246 -2736 2886 -2498
<< via1 >>
rect 1128 -580 1182 -214
rect 1650 -576 1706 -228
rect 1112 -1528 1168 -1374
rect 1646 -1532 1698 -1360
rect 456 -1962 518 -1902
rect 2574 -1896 2626 -1886
rect 2568 -1954 2626 -1896
rect 2574 -1964 2626 -1954
<< metal2 >>
rect 1120 -196 1182 -194
rect 1097 -214 1182 -196
rect 1097 -580 1128 -214
rect 1097 -596 1182 -580
rect 1646 -228 1710 -212
rect 1646 -576 1650 -228
rect 1706 -576 1710 -228
rect 1646 -582 1710 -576
rect 1097 -916 1173 -596
rect 1650 -866 1706 -582
rect 746 -1006 1173 -916
rect 1652 -924 1704 -866
rect 746 -1116 1172 -1006
rect 1098 -1374 1172 -1116
rect 1652 -1124 2074 -924
rect 1652 -1344 1704 -1124
rect 1098 -1528 1112 -1374
rect 1168 -1528 1172 -1374
rect 1098 -1542 1172 -1528
rect 1634 -1360 1704 -1344
rect 1634 -1532 1646 -1360
rect 1698 -1532 1704 -1360
rect 1634 -1546 1704 -1532
rect 1652 -1548 1704 -1546
rect 398 -1870 598 -1868
rect 2538 -1870 2690 -1868
rect 398 -1886 2690 -1870
rect 398 -1896 2574 -1886
rect 398 -1902 2568 -1896
rect 398 -1962 456 -1902
rect 518 -1954 2568 -1902
rect 518 -1960 2574 -1954
rect 518 -1962 598 -1960
rect 2538 -1964 2574 -1960
rect 2626 -1964 2690 -1886
rect 2538 -1966 2690 -1964
use sky130_fd_pr__nfet_01v8_6SJULU  XM1
timestamp 1740557227
transform 0 1 1538 1 0 -2237
box -211 -1210 211 1210
use sky130_fd_pr__pfet_01v8_XLV5ZZ  XM2
timestamp 1740557227
transform 1 0 1255 0 1 -395
box -211 -419 211 419
use sky130_fd_pr__pfet_01v8_XLV5ZZ  XM3
timestamp 1740557227
transform 1 0 1571 0 1 -395
box -211 -419 211 419
use sky130_fd_pr__nfet_01v8_V8CAV6  XM4
timestamp 1740557227
transform 1 0 1245 0 1 -1448
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_V8CAV6  XM5
timestamp 1740557227
transform 1 0 1561 0 1 -1448
box -211 -310 211 310
<< labels >>
flabel metal1 1878 -1548 2078 -1348 0 FreeSans 256 180 0 0 vin2
port 5 nsew
flabel metal1 1324 184 1524 384 0 FreeSans 256 180 0 0 VDD
port 0 nsew
flabel metal1 298 -2712 498 -2512 0 FreeSans 256 180 0 0 GND
port 7 nsew
flabel metal1 732 -1566 932 -1366 0 FreeSans 256 180 0 0 vin1
port 4 nsew
rlabel metal2 746 -1116 946 -916 1 vout1
port 2 n
rlabel metal2 1652 -1124 2074 -924 1 vout2
port 3 n
rlabel metal2 398 -1962 456 -1868 1 Vb
port 6 n
rlabel metal1 1318 -2216 1490 -1638 1 virtual_gnd
<< end >>
