magic
tech sky130A
magscale 1 2
timestamp 1740557227
<< error_p >>
rect -29 1072 29 1078
rect -29 1038 -17 1072
rect -29 1032 29 1038
rect -29 -1038 29 -1032
rect -29 -1072 -17 -1038
rect -29 -1078 29 -1072
<< pwell >>
rect -211 -1210 211 1210
<< nmos >>
rect -15 -1000 15 1000
<< ndiff >>
rect -73 988 -15 1000
rect -73 -988 -61 988
rect -27 -988 -15 988
rect -73 -1000 -15 -988
rect 15 988 73 1000
rect 15 -988 27 988
rect 61 -988 73 988
rect 15 -1000 73 -988
<< ndiffc >>
rect -61 -988 -27 988
rect 27 -988 61 988
<< psubdiff >>
rect -175 1140 -79 1174
rect 79 1140 175 1174
rect -175 1078 -141 1140
rect 141 1078 175 1140
rect -175 -1140 -141 -1078
rect 141 -1140 175 -1078
rect -175 -1174 -79 -1140
rect 79 -1174 175 -1140
<< psubdiffcont >>
rect -79 1140 79 1174
rect -175 -1078 -141 1078
rect 141 -1078 175 1078
rect -79 -1174 79 -1140
<< poly >>
rect -33 1072 33 1088
rect -33 1038 -17 1072
rect 17 1038 33 1072
rect -33 1022 33 1038
rect -15 1000 15 1022
rect -15 -1022 15 -1000
rect -33 -1038 33 -1022
rect -33 -1072 -17 -1038
rect 17 -1072 33 -1038
rect -33 -1088 33 -1072
<< polycont >>
rect -17 1038 17 1072
rect -17 -1072 17 -1038
<< locali >>
rect -175 1140 -79 1174
rect 79 1140 175 1174
rect -175 1078 -141 1140
rect 141 1078 175 1140
rect -33 1038 -17 1072
rect 17 1038 33 1072
rect -61 988 -27 1004
rect -61 -1004 -27 -988
rect 27 988 61 1004
rect 27 -1004 61 -988
rect -33 -1072 -17 -1038
rect 17 -1072 33 -1038
rect -175 -1140 -141 -1078
rect 141 -1140 175 -1078
rect -175 -1174 -79 -1140
rect 79 -1174 175 -1140
<< viali >>
rect -17 1038 17 1072
rect -61 -988 -27 988
rect 27 -988 61 988
rect -17 -1072 17 -1038
<< metal1 >>
rect -29 1072 29 1078
rect -29 1038 -17 1072
rect 17 1038 29 1072
rect -29 1032 29 1038
rect -67 988 -21 1000
rect -67 -988 -61 988
rect -27 -988 -21 988
rect -67 -1000 -21 -988
rect 21 988 67 1000
rect 21 -988 27 988
rect 61 -988 67 988
rect 21 -1000 67 -988
rect -29 -1038 29 -1032
rect -29 -1072 -17 -1038
rect 17 -1072 29 -1038
rect -29 -1078 29 -1072
<< properties >>
string FIXED_BBOX -158 -1157 158 1157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
